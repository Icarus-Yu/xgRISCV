// ----------------------------------------------------------------
// instruction_memory.v
//
// 行为级指令存储器（ROM）模型，用于仿真。
// 它会从一个外部文本文件中读取32位的十六进制指令。
// ----------------------------------------------------------------
module instruction_memory (
    input  [6:0] addr,    // 输入：7位地址，可以寻址 2^7 = 128 条指令
    output reg [31:0] dout // 输出：32位指令数据
);

    // 定义一个存储器数组来存放指令。
    // 大小为128个条目，每个条目32位宽。
    // 这个大小与您Vivado IP核中设置的深度(Depth)128相匹配。
    reg [31:0] mem[0:127];

    // --- 初始化模块 ---
    // initial块中的代码在仿真开始时仅执行一次。
    initial begin
        // 使用Verilog的系统任务$readmemh来从文件中读取十六进制数据。
        // 文件名 "instructions.txt" 应该与您存放机器码的文件名完全一致。
        // 该文件需要放在仿真运行的根目录下。
        $readmemh("instructions.txt", mem);
    end

    // --- 读操作 ---
    // 这是一个组合逻辑块，它会持续地根据输入的地址，从存储器中读取数据。
    // 行为上模拟了一个理想的、无延迟的只读存储器。
    always @(*) begin
        dout = mem[addr];
    end

endmodule
